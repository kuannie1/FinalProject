`include "process.v"

/*
	Convert the input coordinates into pixels
	input: an array with coordinate values
	output: 
		pixels?
*/ 

module rasterize();


endmodule